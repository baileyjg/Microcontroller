`timescale 1ns/10ps

module instructionDecoder();

endmodule